module decoder_top
  (
   input wire clk,
   input wire reset
   );
endmodule   
